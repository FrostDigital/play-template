# 2011-12-02 - Heroku does not seem to like space to much, hence the condense format
# 
# Common stuff
#
email=E-mail
username=E-mail
edit=Edit
delete= Delete
password=Password
confirmPassword=Confirm password
passwords.no-match=Passwords does not match
role=Role
save=Save
show-all=Show all
                         

#
# Password reset
#
passwordReset=Reset password
passwordReset.forgot-it=Forgot your password?
passwordReset.info=Please enter your e-mail in order for us to send further details on how you reset your password. 
passwordReset.sent=Further instructions was sent to your e-mail, please check your inbox. Note that it can take up to 5 minutes for mail to arrive.
passwordReset.mail.subject=Instructions to reset your password
passwordReset.mail.body=Visit this URL to reset your password: \nhttp://localhost:9000/password-reset/%s
passwordReset.notFound=Cannot find any user with e-mail address '%s'
passwordReset.reset.success=OK! Your password has been updated. Please login with new password below.
passwordReset.reset.fail=Could not reset password, please make sure that passwords are valid.
passwordReset.na=Password reset does not exist or is not valid


#
# User settings & administration
#
user.create=Add user
user.delete.self=Cannot delete yourself
user.delete.success=User %s was removed
user.save.success=Saved user %s
user.invited=An invitation has been sent to %s
user.invite=Invite user
user.invite.already-exists=User with e-mail already exists 
user.invite.info=Fill in e-mail and role of user. An invitation will be sent to the users e-mail address.


# 
# Invitation
#
invitation=User invitation
invitation.info=Please complete the form below in order to activate your account.
invitation.mail.subject=You have been invited to "My app name here"
invitation.mail.body=Visit this URL to register your account: \nhttp://localhost:9000/invitation/%s
invitation.success=You are now registered, please login with e-mail and password
invitation.fail=Could not complete invitation.